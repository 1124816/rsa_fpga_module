`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/24/2020 03:36:25 PM
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Selector#(parameter RSA_WIDTH = 128, C_S_AXI_DATA_WIDTH = 32)(
    // Axi4Lite Bus
    input  [C_S_AXI_DATA_WIDTH-1:0] SELECT_IN,
    output [RSA_WIDTH-1 : 0] M_OUT,
    output [RSA_WIDTH-1 : 0] E_OUT,
    output [RSA_WIDTH-1 : 0] N_OUT
);

reg M_OUT;
reg E_OUT = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
reg N_OUT = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000;


always @ (SELECT_IN)begin
    case (SELECT_IN)
        32'b11  : M_OUT <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010001010010100000;
        32'b10  : M_OUT <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000100000;
        32'b01  : M_OUT <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000;
        32'b00  : M_OUT <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000;
        default : M_OUT <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000;
  endcase
end
endmodule
